magic
tech scmos
timestamp 1603947136
<< nwell >>
rect 0 14 38 50
rect -12 -9 38 14
rect -1 -94 27 -73
rect -9 -164 38 -148
rect -8 -178 38 -164
<< pwell >>
rect -12 -55 38 -9
rect -1 -128 27 -94
rect -8 -196 38 -178
<< poly >>
rect 10 61 16 63
rect 10 59 12 61
rect 14 59 16 61
rect 7 57 19 59
rect 7 50 9 57
rect 17 50 19 57
rect 7 42 9 44
rect 17 42 19 44
rect 7 40 19 42
rect 12 38 14 40
rect 12 28 14 32
rect 7 14 9 18
rect 17 14 19 18
rect 7 -11 9 1
rect 17 -1 19 1
rect 13 -3 19 -1
rect 13 -5 15 -3
rect 17 -5 19 -3
rect 13 -7 19 -5
rect 7 -13 13 -11
rect 7 -15 9 -13
rect 11 -15 13 -13
rect 7 -17 13 -15
rect -5 -21 -3 -17
rect 7 -21 9 -17
rect 17 -21 19 -7
rect 29 -21 31 -17
rect -5 -64 -3 -41
rect 7 -59 9 -55
rect 17 -59 19 -55
rect 29 -64 31 -41
rect -5 -66 31 -64
rect 10 -68 12 -66
rect 14 -68 16 -66
rect 10 -70 16 -68
rect 7 -78 9 -74
rect 17 -78 19 -74
rect 7 -96 9 -84
rect 17 -86 19 -84
rect 13 -88 19 -86
rect 13 -90 15 -88
rect 17 -90 19 -88
rect 13 -92 19 -90
rect 7 -98 13 -96
rect 7 -100 9 -98
rect 11 -100 13 -98
rect 7 -102 13 -100
rect 7 -104 9 -102
rect 17 -104 19 -92
rect 7 -114 9 -110
rect 17 -114 19 -110
rect 2 -120 19 -118
rect 2 -122 4 -120
rect 6 -122 8 -120
rect 17 -122 19 -120
rect 2 -124 8 -122
rect 17 -132 19 -128
rect -2 -138 4 -136
rect -2 -140 0 -138
rect 2 -140 31 -138
rect -2 -142 4 -140
rect -2 -148 0 -142
rect 8 -148 10 -144
rect 19 -148 21 -144
rect 29 -148 31 -140
rect -2 -158 0 -154
rect 8 -156 10 -154
rect 19 -156 21 -154
rect 6 -158 12 -156
rect 6 -160 8 -158
rect 10 -160 12 -158
rect 6 -162 12 -160
rect 16 -158 22 -156
rect 29 -158 31 -154
rect 16 -160 18 -158
rect 20 -160 22 -158
rect 16 -162 22 -160
rect 8 -166 10 -162
rect 8 -184 10 -172
rect 8 -194 10 -190
<< ndif >>
rect -12 -23 -5 -21
rect -12 -25 -10 -23
rect -8 -25 -5 -23
rect -12 -30 -5 -25
rect -12 -32 -10 -30
rect -8 -32 -5 -30
rect -12 -37 -5 -32
rect -12 -39 -10 -37
rect -8 -39 -5 -37
rect -12 -41 -5 -39
rect -3 -23 7 -21
rect -3 -25 1 -23
rect 3 -25 7 -23
rect -3 -30 7 -25
rect -3 -32 1 -30
rect 3 -32 7 -30
rect -3 -37 7 -32
rect -3 -39 1 -37
rect 3 -39 7 -37
rect -3 -41 7 -39
rect -1 -44 7 -41
rect -1 -46 1 -44
rect 3 -46 7 -44
rect -1 -51 7 -46
rect -1 -53 1 -51
rect 3 -53 7 -51
rect -1 -55 7 -53
rect 9 -23 17 -21
rect 9 -25 12 -23
rect 14 -25 17 -23
rect 9 -30 17 -25
rect 9 -32 12 -30
rect 14 -32 17 -30
rect 9 -37 17 -32
rect 9 -39 12 -37
rect 14 -39 17 -37
rect 9 -44 17 -39
rect 9 -46 12 -44
rect 14 -46 17 -44
rect 9 -51 17 -46
rect 9 -53 12 -51
rect 14 -53 17 -51
rect 9 -55 17 -53
rect 19 -23 29 -21
rect 19 -25 23 -23
rect 25 -25 29 -23
rect 19 -30 29 -25
rect 19 -32 23 -30
rect 25 -32 29 -30
rect 19 -37 29 -32
rect 19 -39 23 -37
rect 25 -39 29 -37
rect 19 -41 29 -39
rect 31 -23 38 -21
rect 31 -25 34 -23
rect 36 -25 38 -23
rect 31 -30 38 -25
rect 31 -32 34 -30
rect 36 -32 38 -30
rect 31 -37 38 -32
rect 31 -39 34 -37
rect 36 -39 38 -37
rect 31 -41 38 -39
rect 19 -44 27 -41
rect 19 -46 23 -44
rect 25 -46 27 -44
rect 19 -51 27 -46
rect 19 -53 23 -51
rect 25 -53 27 -51
rect 19 -55 27 -53
rect -1 -106 7 -104
rect -1 -108 1 -106
rect 3 -108 7 -106
rect -1 -110 7 -108
rect 9 -106 17 -104
rect 9 -108 12 -106
rect 14 -108 17 -106
rect 9 -110 17 -108
rect 19 -106 27 -104
rect 19 -108 23 -106
rect 25 -108 27 -106
rect 19 -110 27 -108
rect 10 -124 17 -122
rect 10 -126 12 -124
rect 14 -126 17 -124
rect 10 -128 17 -126
rect 19 -124 26 -122
rect 19 -126 22 -124
rect 24 -126 26 -124
rect 19 -128 26 -126
rect 1 -186 8 -184
rect 1 -188 3 -186
rect 5 -188 8 -186
rect 1 -190 8 -188
rect 10 -186 17 -184
rect 10 -188 13 -186
rect 15 -188 17 -186
rect 10 -190 17 -188
<< pdif >>
rect 0 48 7 50
rect 0 46 2 48
rect 4 46 7 48
rect 0 44 7 46
rect 9 48 17 50
rect 9 46 12 48
rect 14 46 17 48
rect 9 44 17 46
rect 19 48 26 50
rect 19 46 22 48
rect 24 46 26 48
rect 19 44 26 46
rect 5 36 12 38
rect 5 34 7 36
rect 9 34 12 36
rect 5 32 12 34
rect 14 36 21 38
rect 14 34 17 36
rect 19 34 21 36
rect 14 32 21 34
rect -1 12 7 14
rect -1 10 1 12
rect 3 10 7 12
rect -1 5 7 10
rect -1 3 1 5
rect 3 3 7 5
rect -1 1 7 3
rect 9 12 17 14
rect 9 10 12 12
rect 14 10 17 12
rect 9 5 17 10
rect 9 3 12 5
rect 14 3 17 5
rect 9 1 17 3
rect 19 12 27 14
rect 19 10 23 12
rect 25 10 27 12
rect 19 5 27 10
rect 19 3 23 5
rect 25 3 27 5
rect 19 1 27 3
rect -1 -80 7 -78
rect -1 -82 1 -80
rect 3 -82 7 -80
rect -1 -84 7 -82
rect 9 -80 17 -78
rect 9 -82 12 -80
rect 14 -82 17 -80
rect 9 -84 17 -82
rect 19 -80 27 -78
rect 19 -82 23 -80
rect 25 -82 27 -80
rect 19 -84 27 -82
rect -9 -150 -2 -148
rect -9 -152 -7 -150
rect -5 -152 -2 -150
rect -9 -154 -2 -152
rect 0 -150 8 -148
rect 0 -152 3 -150
rect 5 -152 8 -150
rect 0 -154 8 -152
rect 10 -150 19 -148
rect 10 -152 14 -150
rect 16 -152 19 -150
rect 10 -154 19 -152
rect 21 -150 29 -148
rect 21 -152 24 -150
rect 26 -152 29 -150
rect 21 -154 29 -152
rect 31 -150 38 -148
rect 31 -152 34 -150
rect 36 -152 38 -150
rect 31 -154 38 -152
rect 1 -168 8 -166
rect 1 -170 3 -168
rect 5 -170 8 -168
rect 1 -172 8 -170
rect 10 -168 17 -166
rect 10 -170 13 -168
rect 15 -170 17 -168
rect 10 -172 17 -170
<< alu1 >>
rect 11 61 15 62
rect 11 59 12 61
rect 14 59 15 61
rect 11 58 15 59
rect 11 53 15 54
rect 11 51 12 53
rect 14 51 15 53
rect 1 48 5 49
rect 1 46 2 48
rect 4 46 5 48
rect 1 37 5 46
rect 11 48 15 51
rect 11 46 12 48
rect 14 46 15 48
rect 11 45 15 46
rect 21 48 25 49
rect 21 46 22 48
rect 24 46 25 48
rect 21 37 25 46
rect -11 36 10 37
rect -11 34 7 36
rect 9 34 10 36
rect -11 33 10 34
rect 16 36 37 37
rect 16 34 17 36
rect 19 34 37 36
rect 16 33 37 34
rect -11 -23 -7 33
rect 11 19 15 20
rect 11 17 12 19
rect 14 17 15 19
rect -11 -25 -10 -23
rect -8 -25 -7 -23
rect -11 -30 -7 -25
rect -11 -32 -10 -30
rect -8 -32 -7 -30
rect -11 -37 -7 -32
rect -11 -39 -10 -37
rect -8 -39 -7 -37
rect -11 -97 -7 -39
rect 0 12 4 13
rect 0 10 1 12
rect 3 10 4 12
rect 0 5 4 10
rect 0 3 1 5
rect 3 3 4 5
rect 0 -2 4 3
rect 11 12 15 17
rect 11 10 12 12
rect 14 10 15 12
rect 11 5 15 10
rect 11 3 12 5
rect 14 3 15 5
rect 11 2 15 3
rect 22 12 26 13
rect 22 10 23 12
rect 25 10 26 12
rect 22 5 26 10
rect 22 3 23 5
rect 25 3 26 5
rect 0 -3 18 -2
rect 0 -5 15 -3
rect 17 -5 18 -3
rect 0 -6 18 -5
rect 0 -23 4 -6
rect 22 -12 26 3
rect 8 -13 26 -12
rect 8 -15 9 -13
rect 11 -15 26 -13
rect 8 -16 26 -15
rect 0 -25 1 -23
rect 3 -25 4 -23
rect 0 -30 4 -25
rect 0 -32 1 -30
rect 3 -32 4 -30
rect 0 -37 4 -32
rect 0 -39 1 -37
rect 3 -39 4 -37
rect 0 -44 4 -39
rect 0 -46 1 -44
rect 3 -46 4 -44
rect 0 -51 4 -46
rect 0 -53 1 -51
rect 3 -53 4 -51
rect 0 -54 4 -53
rect 11 -23 15 -22
rect 11 -25 12 -23
rect 14 -25 15 -23
rect 11 -30 15 -25
rect 11 -32 12 -30
rect 14 -32 15 -30
rect 11 -37 15 -32
rect 11 -39 12 -37
rect 14 -39 15 -37
rect 11 -44 15 -39
rect 11 -46 12 -44
rect 14 -46 15 -44
rect 11 -51 15 -46
rect 11 -53 12 -51
rect 14 -53 15 -51
rect 11 -58 15 -53
rect 22 -23 26 -16
rect 22 -25 23 -23
rect 25 -25 26 -23
rect 22 -30 26 -25
rect 22 -32 23 -30
rect 25 -32 26 -30
rect 22 -37 26 -32
rect 22 -39 23 -37
rect 25 -39 26 -37
rect 22 -44 26 -39
rect 22 -46 23 -44
rect 25 -46 26 -44
rect 22 -51 26 -46
rect 22 -53 23 -51
rect 25 -53 26 -51
rect 22 -54 26 -53
rect 33 -23 37 33
rect 33 -25 34 -23
rect 36 -25 37 -23
rect 33 -30 37 -25
rect 33 -32 34 -30
rect 36 -32 37 -30
rect 33 -37 37 -32
rect 33 -39 34 -37
rect 36 -39 37 -37
rect 11 -60 12 -58
rect 14 -60 15 -58
rect 11 -61 15 -60
rect 11 -66 15 -65
rect 11 -68 12 -66
rect 14 -68 15 -66
rect 11 -69 15 -68
rect 11 -74 15 -73
rect 11 -76 12 -74
rect 14 -76 15 -74
rect 0 -80 4 -79
rect 0 -82 1 -80
rect 3 -82 4 -80
rect 0 -87 4 -82
rect 11 -80 15 -76
rect 11 -82 12 -80
rect 14 -82 15 -80
rect 11 -83 15 -82
rect 22 -80 26 -79
rect 22 -82 23 -80
rect 25 -82 26 -80
rect 22 -87 26 -82
rect 33 -87 37 -39
rect 0 -88 18 -87
rect 0 -90 15 -88
rect 17 -90 18 -88
rect 0 -91 18 -90
rect 22 -91 37 -87
rect 0 -97 4 -91
rect 22 -97 26 -91
rect -11 -101 4 -97
rect 8 -98 26 -97
rect 8 -100 9 -98
rect 11 -100 26 -98
rect 8 -101 26 -100
rect -11 -149 -7 -101
rect 0 -106 4 -101
rect 0 -108 1 -106
rect 3 -108 4 -106
rect 0 -109 4 -108
rect 11 -106 15 -105
rect 11 -108 12 -106
rect 14 -108 15 -106
rect 3 -120 7 -119
rect 3 -122 4 -120
rect 6 -122 7 -120
rect 3 -123 7 -122
rect 11 -124 15 -108
rect 22 -106 26 -101
rect 22 -108 23 -106
rect 25 -108 26 -106
rect 22 -109 26 -108
rect 11 -126 12 -124
rect 14 -126 15 -124
rect 11 -127 15 -126
rect 21 -124 25 -123
rect 21 -126 22 -124
rect 24 -126 25 -124
rect 21 -129 25 -126
rect 21 -131 22 -129
rect 24 -131 25 -129
rect 21 -132 25 -131
rect -1 -138 3 -137
rect -1 -140 0 -138
rect 2 -140 3 -138
rect -1 -141 3 -140
rect -11 -150 -4 -149
rect -11 -152 -7 -150
rect -5 -152 -4 -150
rect -11 -153 -4 -152
rect 2 -150 6 -149
rect 2 -152 3 -150
rect 5 -152 6 -150
rect 2 -153 6 -152
rect 13 -150 17 -149
rect 13 -152 14 -150
rect 16 -152 17 -150
rect 13 -153 17 -152
rect 23 -150 27 -149
rect 23 -152 24 -150
rect 26 -152 27 -150
rect 23 -153 27 -152
rect 33 -150 37 -91
rect 33 -152 34 -150
rect 36 -152 37 -150
rect -11 -196 -7 -153
rect 7 -158 11 -157
rect 7 -160 8 -158
rect 10 -160 11 -158
rect 7 -161 11 -160
rect 17 -158 21 -157
rect 17 -160 18 -158
rect 20 -160 21 -158
rect 17 -167 21 -160
rect 2 -168 6 -167
rect 2 -170 3 -168
rect 5 -170 6 -168
rect 2 -171 6 -170
rect 12 -168 21 -167
rect 12 -170 13 -168
rect 15 -170 21 -168
rect 12 -171 21 -170
rect 25 -160 29 -159
rect 25 -162 26 -160
rect 28 -162 29 -160
rect 2 -186 6 -185
rect 2 -188 3 -186
rect 5 -188 6 -186
rect 2 -189 6 -188
rect 12 -186 16 -171
rect 12 -188 13 -186
rect 15 -188 16 -186
rect 12 -189 16 -188
rect 25 -186 29 -162
rect 25 -188 26 -186
rect 28 -188 29 -186
rect 25 -189 29 -188
rect 33 -196 37 -152
<< alu2 >>
rect -11 61 37 62
rect -11 59 12 61
rect 14 59 37 61
rect -11 58 37 59
rect -23 53 41 54
rect -23 51 12 53
rect 14 51 41 53
rect -23 50 41 51
rect -23 20 -19 50
rect -23 19 41 20
rect -23 17 12 19
rect 14 17 41 19
rect -23 16 41 17
rect -23 -73 -19 16
rect 45 -57 49 50
rect -15 -58 49 -57
rect -15 -60 12 -58
rect 14 -60 49 -58
rect -15 -61 49 -60
rect -15 -66 41 -65
rect -15 -68 12 -66
rect 14 -68 41 -66
rect -15 -69 41 -68
rect -23 -74 41 -73
rect -23 -76 12 -74
rect 14 -76 41 -74
rect -23 -77 41 -76
rect -23 -167 -19 -77
rect -15 -120 41 -119
rect -15 -122 4 -120
rect 6 -122 41 -120
rect -15 -123 41 -122
rect 45 -128 49 -61
rect -15 -129 49 -128
rect -15 -131 22 -129
rect 24 -131 49 -129
rect -15 -132 49 -131
rect -15 -138 41 -137
rect -15 -140 0 -138
rect 2 -140 41 -138
rect -15 -141 41 -140
rect 13 -150 29 -149
rect 13 -152 14 -150
rect 16 -152 29 -150
rect 13 -153 29 -152
rect -15 -158 11 -157
rect -15 -160 8 -158
rect 10 -160 11 -158
rect -15 -161 11 -160
rect 25 -160 29 -153
rect 25 -162 26 -160
rect 28 -162 29 -160
rect 25 -163 29 -162
rect -23 -168 6 -167
rect -23 -170 3 -168
rect 5 -170 6 -168
rect -23 -171 6 -170
rect -23 -189 -19 -171
rect 2 -172 6 -171
rect 21 -171 41 -167
rect 21 -172 25 -171
rect 2 -176 25 -172
rect 2 -184 25 -180
rect 2 -185 6 -184
rect -15 -186 6 -185
rect -15 -188 3 -186
rect 5 -188 6 -186
rect -15 -189 6 -188
rect 21 -185 25 -184
rect 45 -185 49 -132
rect 21 -186 49 -185
rect 21 -188 26 -186
rect 28 -188 49 -186
rect 21 -189 49 -188
<< nmos >>
rect -5 -41 -3 -21
rect 7 -55 9 -21
rect 17 -55 19 -21
rect 29 -41 31 -21
rect 7 -110 9 -104
rect 17 -110 19 -104
rect 17 -128 19 -122
rect 8 -190 10 -184
<< pmos >>
rect 7 44 9 50
rect 17 44 19 50
rect 12 32 14 38
rect 7 1 9 14
rect 17 1 19 14
rect 7 -84 9 -78
rect 17 -84 19 -78
rect -2 -154 0 -148
rect 8 -154 10 -148
rect 19 -154 21 -148
rect 29 -154 31 -148
rect 8 -172 10 -166
<< polyct1 >>
rect 12 59 14 61
rect 15 -5 17 -3
rect 9 -15 11 -13
rect 12 -68 14 -66
rect 15 -90 17 -88
rect 9 -100 11 -98
rect 4 -122 6 -120
rect 0 -140 2 -138
rect 8 -160 10 -158
rect 18 -160 20 -158
<< ndifct1 >>
rect -10 -25 -8 -23
rect -10 -32 -8 -30
rect -10 -39 -8 -37
rect 1 -25 3 -23
rect 1 -32 3 -30
rect 1 -39 3 -37
rect 1 -46 3 -44
rect 1 -53 3 -51
rect 12 -25 14 -23
rect 12 -32 14 -30
rect 12 -39 14 -37
rect 12 -46 14 -44
rect 12 -53 14 -51
rect 23 -25 25 -23
rect 23 -32 25 -30
rect 23 -39 25 -37
rect 34 -25 36 -23
rect 34 -32 36 -30
rect 34 -39 36 -37
rect 23 -46 25 -44
rect 23 -53 25 -51
rect 1 -108 3 -106
rect 12 -108 14 -106
rect 23 -108 25 -106
rect 12 -126 14 -124
rect 22 -126 24 -124
rect 3 -188 5 -186
rect 13 -188 15 -186
<< pdifct1 >>
rect 2 46 4 48
rect 12 46 14 48
rect 22 46 24 48
rect 7 34 9 36
rect 17 34 19 36
rect 1 10 3 12
rect 1 3 3 5
rect 12 10 14 12
rect 12 3 14 5
rect 23 10 25 12
rect 23 3 25 5
rect 1 -82 3 -80
rect 12 -82 14 -80
rect 23 -82 25 -80
rect -7 -152 -5 -150
rect 3 -152 5 -150
rect 14 -152 16 -150
rect 24 -152 26 -150
rect 34 -152 36 -150
rect 3 -170 5 -168
rect 13 -170 15 -168
<< via1 >>
rect 12 59 14 61
rect 12 51 14 53
rect 12 17 14 19
rect 12 -60 14 -58
rect 12 -68 14 -66
rect 12 -76 14 -74
rect 4 -122 6 -120
rect 22 -131 24 -129
rect 0 -140 2 -138
rect 14 -152 16 -150
rect 8 -160 10 -158
rect 3 -170 5 -168
rect 26 -162 28 -160
rect 3 -188 5 -186
rect 26 -188 28 -186
<< labels >>
rlabel alu1 -9 22 -9 22 5 BL
rlabel alu1 35 22 35 22 5 BLB
rlabel via1 13 18 13 18 1 Vdd
rlabel via1 13 -59 13 -59 1 Gnd
rlabel via1 13 -67 13 -67 1 WL
rlabel via1 5 -121 5 -121 1 SAE
rlabel via1 23 -130 23 -130 1 Gnd
rlabel via1 13 -75 13 -75 1 Vdd
rlabel alu1 -9 -71 -9 -71 5 BL
rlabel alu1 35 -71 35 -71 5 BLB
rlabel via1 4 -169 4 -169 1 Vdd
rlabel via1 4 -187 4 -187 1 Gnd
rlabel via1 1 -139 1 -139 1 WE
rlabel alu1 -9 -134 -9 -134 5 BL
rlabel alu1 35 -134 35 -134 5 BLB
rlabel alu1 -9 -191 -9 -191 1 BL
rlabel alu1 35 -191 35 -191 1 BLB
rlabel via1 9 -159 9 -159 1 DATA
rlabel alu1 2 -4 2 -4 1 A
rlabel alu1 24 -4 24 -4 1 AB
rlabel alu1 -9 35 -9 35 3 BL
rlabel alu1 35 35 35 35 7 BLB
rlabel via1 13 52 13 52 1 Vdd
rlabel via1 13 60 13 60 5 PRE
<< end >>
