magic
tech scmos
timestamp 1603894115
<< nwell >>
rect -13 -1 13 17
<< poly >>
rect -3 28 3 30
rect -3 26 -1 28
rect 1 26 3 28
rect -6 24 6 26
rect -6 17 -4 24
rect 4 17 6 24
rect -6 9 -4 11
rect 4 9 6 11
rect -6 7 6 9
rect -1 5 1 7
rect -1 -5 1 -1
<< pdif >>
rect -13 15 -6 17
rect -13 13 -11 15
rect -9 13 -6 15
rect -13 11 -6 13
rect -4 15 4 17
rect -4 13 -1 15
rect 1 13 4 15
rect -4 11 4 13
rect 6 15 13 17
rect 6 13 9 15
rect 11 13 13 15
rect 6 11 13 13
rect -8 3 -1 5
rect -8 1 -6 3
rect -4 1 -1 3
rect -8 -1 -1 1
rect 1 3 8 5
rect 1 1 4 3
rect 6 1 8 3
rect 1 -1 8 1
<< alu1 >>
rect -2 28 2 29
rect -2 26 -1 28
rect 1 26 2 28
rect -2 25 2 26
rect -2 20 2 21
rect -2 18 -1 20
rect 1 18 2 20
rect -12 15 -8 16
rect -12 13 -11 15
rect -9 13 -8 15
rect -12 4 -8 13
rect -2 15 2 18
rect -2 13 -1 15
rect 1 13 2 15
rect -2 12 2 13
rect 8 15 12 16
rect 8 13 9 15
rect 11 13 12 15
rect 8 4 12 13
rect -24 3 -3 4
rect -24 1 -6 3
rect -4 1 -3 3
rect -24 0 -3 1
rect 3 3 24 4
rect 3 1 4 3
rect 6 1 24 3
rect 3 0 24 1
rect -24 -8 -20 0
rect 20 -8 24 0
<< alu2 >>
rect -24 28 24 29
rect -24 26 -1 28
rect 1 26 24 28
rect -24 25 24 26
rect -24 20 24 21
rect -24 18 -1 20
rect 1 18 24 20
rect -24 17 24 18
<< pmos >>
rect -6 11 -4 17
rect 4 11 6 17
rect -1 -1 1 5
<< polyct1 >>
rect -1 26 1 28
<< pdifct1 >>
rect -11 13 -9 15
rect -1 13 1 15
rect 9 13 11 15
rect -6 1 -4 3
rect 4 1 6 3
<< via1 >>
rect -1 26 1 28
rect -1 18 1 20
<< labels >>
rlabel alu1 -22 2 -22 2 3 BL
rlabel alu1 22 2 22 2 7 BLB
rlabel via1 0 19 0 19 1 Vdd
rlabel via1 0 27 0 27 5 PRE
<< end >>
