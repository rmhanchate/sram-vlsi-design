magic
tech scmos
timestamp 1603920245
<< nwell >>
rect -35 10 15 33
<< pwell >>
rect -35 -36 15 10
<< poly >>
rect -16 33 -14 37
rect -6 33 -4 37
rect -16 8 -14 20
rect -6 18 -4 20
rect -10 16 -4 18
rect -10 14 -8 16
rect -6 14 -4 16
rect -10 12 -4 14
rect -16 6 -10 8
rect -16 4 -14 6
rect -12 4 -10 6
rect -16 2 -10 4
rect -28 -2 -26 2
rect -16 -2 -14 2
rect -6 -2 -4 12
rect 6 -2 8 2
rect -28 -45 -26 -22
rect -16 -40 -14 -36
rect -6 -40 -4 -36
rect 6 -45 8 -22
rect -28 -47 8 -45
rect -13 -49 -11 -47
rect -9 -49 -7 -47
rect -13 -51 -7 -49
<< ndif >>
rect -35 -4 -28 -2
rect -35 -6 -33 -4
rect -31 -6 -28 -4
rect -35 -11 -28 -6
rect -35 -13 -33 -11
rect -31 -13 -28 -11
rect -35 -18 -28 -13
rect -35 -20 -33 -18
rect -31 -20 -28 -18
rect -35 -22 -28 -20
rect -26 -4 -16 -2
rect -26 -6 -22 -4
rect -20 -6 -16 -4
rect -26 -11 -16 -6
rect -26 -13 -22 -11
rect -20 -13 -16 -11
rect -26 -18 -16 -13
rect -26 -20 -22 -18
rect -20 -20 -16 -18
rect -26 -22 -16 -20
rect -24 -25 -16 -22
rect -24 -27 -22 -25
rect -20 -27 -16 -25
rect -24 -32 -16 -27
rect -24 -34 -22 -32
rect -20 -34 -16 -32
rect -24 -36 -16 -34
rect -14 -4 -6 -2
rect -14 -6 -11 -4
rect -9 -6 -6 -4
rect -14 -11 -6 -6
rect -14 -13 -11 -11
rect -9 -13 -6 -11
rect -14 -18 -6 -13
rect -14 -20 -11 -18
rect -9 -20 -6 -18
rect -14 -25 -6 -20
rect -14 -27 -11 -25
rect -9 -27 -6 -25
rect -14 -32 -6 -27
rect -14 -34 -11 -32
rect -9 -34 -6 -32
rect -14 -36 -6 -34
rect -4 -4 6 -2
rect -4 -6 0 -4
rect 2 -6 6 -4
rect -4 -11 6 -6
rect -4 -13 0 -11
rect 2 -13 6 -11
rect -4 -18 6 -13
rect -4 -20 0 -18
rect 2 -20 6 -18
rect -4 -22 6 -20
rect 8 -4 15 -2
rect 8 -6 11 -4
rect 13 -6 15 -4
rect 8 -11 15 -6
rect 8 -13 11 -11
rect 13 -13 15 -11
rect 8 -18 15 -13
rect 8 -20 11 -18
rect 13 -20 15 -18
rect 8 -22 15 -20
rect -4 -25 4 -22
rect -4 -27 0 -25
rect 2 -27 4 -25
rect -4 -32 4 -27
rect -4 -34 0 -32
rect 2 -34 4 -32
rect -4 -36 4 -34
<< pdif >>
rect -24 31 -16 33
rect -24 29 -22 31
rect -20 29 -16 31
rect -24 24 -16 29
rect -24 22 -22 24
rect -20 22 -16 24
rect -24 20 -16 22
rect -14 31 -6 33
rect -14 29 -11 31
rect -9 29 -6 31
rect -14 24 -6 29
rect -14 22 -11 24
rect -9 22 -6 24
rect -14 20 -6 22
rect -4 31 4 33
rect -4 29 0 31
rect 2 29 4 31
rect -4 24 4 29
rect -4 22 0 24
rect 2 22 4 24
rect -4 20 4 22
<< alu1 >>
rect -34 -4 -30 43
rect -12 38 -8 39
rect -12 36 -11 38
rect -9 36 -8 38
rect -34 -6 -33 -4
rect -31 -6 -30 -4
rect -34 -11 -30 -6
rect -34 -13 -33 -11
rect -31 -13 -30 -11
rect -34 -18 -30 -13
rect -34 -20 -33 -18
rect -31 -20 -30 -18
rect -34 -54 -30 -20
rect -23 31 -19 32
rect -23 29 -22 31
rect -20 29 -19 31
rect -23 24 -19 29
rect -23 22 -22 24
rect -20 22 -19 24
rect -23 17 -19 22
rect -12 31 -8 36
rect -12 29 -11 31
rect -9 29 -8 31
rect -12 24 -8 29
rect -12 22 -11 24
rect -9 22 -8 24
rect -12 21 -8 22
rect -1 31 3 32
rect -1 29 0 31
rect 2 29 3 31
rect -1 24 3 29
rect -1 22 0 24
rect 2 22 3 24
rect -23 16 -5 17
rect -23 14 -8 16
rect -6 14 -5 16
rect -23 13 -5 14
rect -23 -4 -19 13
rect -1 7 3 22
rect -15 6 3 7
rect -15 4 -14 6
rect -12 4 3 6
rect -15 3 3 4
rect -23 -6 -22 -4
rect -20 -6 -19 -4
rect -23 -11 -19 -6
rect -23 -13 -22 -11
rect -20 -13 -19 -11
rect -23 -18 -19 -13
rect -23 -20 -22 -18
rect -20 -20 -19 -18
rect -23 -25 -19 -20
rect -23 -27 -22 -25
rect -20 -27 -19 -25
rect -23 -32 -19 -27
rect -23 -34 -22 -32
rect -20 -34 -19 -32
rect -23 -35 -19 -34
rect -12 -4 -8 -3
rect -12 -6 -11 -4
rect -9 -6 -8 -4
rect -12 -11 -8 -6
rect -12 -13 -11 -11
rect -9 -13 -8 -11
rect -12 -18 -8 -13
rect -12 -20 -11 -18
rect -9 -20 -8 -18
rect -12 -25 -8 -20
rect -12 -27 -11 -25
rect -9 -27 -8 -25
rect -12 -32 -8 -27
rect -12 -34 -11 -32
rect -9 -34 -8 -32
rect -12 -39 -8 -34
rect -1 -4 3 3
rect -1 -6 0 -4
rect 2 -6 3 -4
rect -1 -11 3 -6
rect -1 -13 0 -11
rect 2 -13 3 -11
rect -1 -18 3 -13
rect -1 -20 0 -18
rect 2 -20 3 -18
rect -1 -25 3 -20
rect -1 -27 0 -25
rect 2 -27 3 -25
rect -1 -32 3 -27
rect -1 -34 0 -32
rect 2 -34 3 -32
rect -1 -35 3 -34
rect 10 -4 14 43
rect 10 -6 11 -4
rect 13 -6 14 -4
rect 10 -11 14 -6
rect 10 -13 11 -11
rect 13 -13 14 -11
rect 10 -18 14 -13
rect 10 -20 11 -18
rect 13 -20 14 -18
rect -12 -41 -11 -39
rect -9 -41 -8 -39
rect -12 -42 -8 -41
rect -12 -47 -8 -46
rect -12 -49 -11 -47
rect -9 -49 -8 -47
rect -12 -50 -8 -49
rect 10 -54 14 -20
<< alu2 >>
rect -38 38 18 39
rect -38 36 -11 38
rect -9 36 18 38
rect -38 35 18 36
rect -38 -39 18 -38
rect -38 -41 -11 -39
rect -9 -41 18 -39
rect -38 -42 18 -41
rect -38 -47 18 -46
rect -38 -49 -11 -47
rect -9 -49 18 -47
rect -38 -50 18 -49
<< nmos >>
rect -28 -22 -26 -2
rect -16 -36 -14 -2
rect -6 -36 -4 -2
rect 6 -22 8 -2
<< pmos >>
rect -16 20 -14 33
rect -6 20 -4 33
<< polyct1 >>
rect -8 14 -6 16
rect -14 4 -12 6
rect -11 -49 -9 -47
<< ndifct1 >>
rect -33 -6 -31 -4
rect -33 -13 -31 -11
rect -33 -20 -31 -18
rect -22 -6 -20 -4
rect -22 -13 -20 -11
rect -22 -20 -20 -18
rect -22 -27 -20 -25
rect -22 -34 -20 -32
rect -11 -6 -9 -4
rect -11 -13 -9 -11
rect -11 -20 -9 -18
rect -11 -27 -9 -25
rect -11 -34 -9 -32
rect 0 -6 2 -4
rect 0 -13 2 -11
rect 0 -20 2 -18
rect 11 -6 13 -4
rect 11 -13 13 -11
rect 11 -20 13 -18
rect 0 -27 2 -25
rect 0 -34 2 -32
<< pdifct1 >>
rect -22 29 -20 31
rect -22 22 -20 24
rect -11 29 -9 31
rect -11 22 -9 24
rect 0 29 2 31
rect 0 22 2 24
<< via1 >>
rect -11 36 -9 38
rect -11 -41 -9 -39
rect -11 -49 -9 -47
<< labels >>
rlabel alu1 -32 41 -32 41 5 BL
rlabel alu1 12 41 12 41 5 BLB
rlabel via1 -10 37 -10 37 1 Vdd
rlabel via1 -10 -40 -10 -40 1 Gnd
rlabel via1 -10 -48 -10 -48 1 WL
rlabel alu1 -32 -52 -32 -52 1 BL
rlabel alu1 12 -52 12 -52 1 BLB
rlabel alu1 -21 15 -21 15 1 A
rlabel alu1 1 15 1 15 1 AB
<< end >>
