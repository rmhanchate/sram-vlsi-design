magic
tech scmos
timestamp 1603896608
<< nwell >>
rect -14 0 14 21
<< pwell >>
rect -14 -34 14 0
<< poly >>
rect -6 16 -4 20
rect 4 16 6 20
rect -6 -2 -4 10
rect 4 8 6 10
rect 0 6 6 8
rect 0 4 2 6
rect 4 4 6 6
rect 0 2 6 4
rect -6 -4 0 -2
rect -6 -6 -4 -4
rect -2 -6 0 -4
rect -6 -8 0 -6
rect -6 -10 -4 -8
rect 4 -10 6 2
rect -6 -20 -4 -16
rect 4 -20 6 -16
rect -11 -26 6 -24
rect -11 -28 -9 -26
rect -7 -28 -5 -26
rect 4 -28 6 -26
rect -11 -30 -5 -28
rect 4 -38 6 -34
<< ndif >>
rect -14 -12 -6 -10
rect -14 -14 -12 -12
rect -10 -14 -6 -12
rect -14 -16 -6 -14
rect -4 -12 4 -10
rect -4 -14 -1 -12
rect 1 -14 4 -12
rect -4 -16 4 -14
rect 6 -12 14 -10
rect 6 -14 10 -12
rect 12 -14 14 -12
rect 6 -16 14 -14
rect -3 -30 4 -28
rect -3 -32 -1 -30
rect 1 -32 4 -30
rect -3 -34 4 -32
rect 6 -30 13 -28
rect 6 -32 9 -30
rect 11 -32 13 -30
rect 6 -34 13 -32
<< pdif >>
rect -14 14 -6 16
rect -14 12 -12 14
rect -10 12 -6 14
rect -14 10 -6 12
rect -4 14 4 16
rect -4 12 -1 14
rect 1 12 4 14
rect -4 10 4 12
rect 6 14 14 16
rect 6 12 10 14
rect 12 12 14 14
rect 6 10 14 12
<< alu1 >>
rect -24 -3 -20 25
rect -2 20 2 21
rect -2 18 -1 20
rect 1 18 2 20
rect -13 14 -9 15
rect -13 12 -12 14
rect -10 12 -9 14
rect -13 7 -9 12
rect -2 14 2 18
rect -2 12 -1 14
rect 1 12 2 14
rect -2 11 2 12
rect 9 14 13 15
rect 9 12 10 14
rect 12 12 13 14
rect 9 7 13 12
rect 20 7 24 25
rect -13 6 5 7
rect -13 4 2 6
rect 4 4 5 6
rect -13 3 5 4
rect 9 3 24 7
rect -13 -3 -9 3
rect 9 -3 13 3
rect -24 -7 -9 -3
rect -5 -4 13 -3
rect -5 -6 -4 -4
rect -2 -6 13 -4
rect -5 -7 13 -6
rect -24 -42 -20 -7
rect -13 -12 -9 -7
rect -13 -14 -12 -12
rect -10 -14 -9 -12
rect -13 -15 -9 -14
rect -2 -12 2 -11
rect -2 -14 -1 -12
rect 1 -14 2 -12
rect -10 -26 -6 -25
rect -10 -28 -9 -26
rect -7 -28 -6 -26
rect -10 -29 -6 -28
rect -2 -30 2 -14
rect 9 -12 13 -7
rect 9 -14 10 -12
rect 12 -14 13 -12
rect 9 -15 13 -14
rect -2 -32 -1 -30
rect 1 -32 2 -30
rect -2 -33 2 -32
rect 8 -30 12 -29
rect 8 -32 9 -30
rect 11 -32 12 -30
rect 8 -35 12 -32
rect 8 -37 9 -35
rect 11 -37 12 -35
rect 8 -38 12 -37
rect 20 -42 24 3
<< alu2 >>
rect -28 20 28 21
rect -28 18 -1 20
rect 1 18 28 20
rect -28 17 28 18
rect -28 -26 28 -25
rect -28 -28 -9 -26
rect -7 -28 28 -26
rect -28 -29 28 -28
rect -28 -35 28 -34
rect -28 -37 9 -35
rect 11 -37 28 -35
rect -28 -38 28 -37
<< nmos >>
rect -6 -16 -4 -10
rect 4 -16 6 -10
rect 4 -34 6 -28
<< pmos >>
rect -6 10 -4 16
rect 4 10 6 16
<< polyct1 >>
rect 2 4 4 6
rect -4 -6 -2 -4
rect -9 -28 -7 -26
<< ndifct1 >>
rect -12 -14 -10 -12
rect -1 -14 1 -12
rect 10 -14 12 -12
rect -1 -32 1 -30
rect 9 -32 11 -30
<< pdifct1 >>
rect -12 12 -10 14
rect -1 12 1 14
rect 10 12 12 14
<< via1 >>
rect -1 18 1 20
rect -9 -28 -7 -26
rect 9 -37 11 -35
<< labels >>
rlabel via1 -8 -27 -8 -27 1 SAE
rlabel via1 10 -36 10 -36 1 Gnd
rlabel via1 0 19 0 19 1 Vdd
rlabel alu1 -22 23 -22 23 5 BL
rlabel alu1 22 23 22 23 5 BLB
rlabel alu1 -22 -40 -22 -40 1 BL
rlabel alu1 22 -40 22 -40 1 BLB
<< end >>
